// https://eprint.iacr.org/2011/332.pdf
// And http://cs-www.cs.yale.edu/homes/peralta/CircuitStuff/AESDEPTH16SIZE125
// But much larger than a simple LUT based approach.

module tiny_sbox
(
    input wire [7:0] in,
    output wire [7:0] out
);

    // 1 bit elements:
    // + corresponds to XOR
    // x corresponds to AND
    // # means XNOR, or ~^

    wire [7:0] x;
    assign x[0] = in[7];
    assign x[1] = in[6];
    assign x[2] = in[5];
    assign x[3] = in[4];
    assign x[4] = in[3];
    assign x[5] = in[2];
    assign x[6] = in[1];
    assign x[7] = in[0];

    // T1 = U6 + U4
    wire T1 = x[6] ^ x[4];
    // T2 = U3 + U0
    wire T2 = x[3] ^ x[0];
    // T3 = U1 + U2
    wire T3 = x[1] ^ x[2];
    // T4 = U7 + T3
    wire T4 = x[7] ^ T3;
    // T5 = T1 + T2
    wire T5 = T1 ^ T2;
    // T6 = U1 + U5
    wire T6 = x[1] ^ x[5];
    // T7 = U0 + U6
    wire T7 = x[0] ^ x[6];
    // T8 = T1 + T6
    wire T8 = T1 ^ T6;
    // T9 = U6 + T4
    wire T9 = x[6] ^ T4;
    // T10 = U3 + T4
    wire T10 = x[3] ^ T4;
    // T11 = U7 + T5
    wire T11 = x[7] ^ T5;
    // T12 = T5 + T6
    wire T12 = T5 ^ T6;
    // T13 = U2 + U5
    wire T13 = x[2] ^ x[5];
    // T14 = T3 + T5
    wire T14 = T3 ^ T5;
    // T15 = U5 + T7
    wire T15 = x[5] ^ T7;
    // T16 = U0 + U5
    wire T16 = x[0] ^ x[5];
    // T17 = U7 + T8
    wire T17 = x[7] ^ T8;
    // T18 = U6 + U5
    wire T18 = x[6] ^ x[5];
    // T19 = T2 + T18
    wire T19 = T2 ^ T18;
    // T20 = T4 + T15
    wire T20 = T4 ^ T15;
    // T21 = T1 + T13
    wire T21 = T1 ^ T13;
    // T22 = U0 + T4
    wire T22 = x[0] ^ T4;
    // T39 = T21 + T5
    wire T39 = T21 ^ T5;
    // T40 = T21 + T7
    wire T40 = T21 ^ T7;
    // T41 = T7 + T19
    wire T41 = T7 ^ T19;
    // T42 = T16 + T14
    wire T42 = T16 ^ T14;
    // T43 = T22 + T17
    wire T43 = T22 ^ T17;
    // T44 = T19 x T5
    wire T44 = T19 & T5;
    // T45 = T20 x T11
    wire T45 = T20 & T11;
    // T46 = T12 + T44
    wire T46 = T12 ^ T44;
    // T47 = T10 x U7
    wire T47 = T10 & x[7];
    // T48 = T47 + T44
    wire T48 = T47 ^ T44;
    // T49 = T7 x T21
    wire T49 = T7 & T21;
    // T50 = T9 x T4
    wire T50 = T9 & T4;
    // T51 = T40 + T49
    wire T51 = T40 ^ T49;
    // T52 = T22 x T17
    wire T52 = T22 & T17;
    // T53 = T52 + T49
    wire T53 = T52 ^ T49;
    // T54 = T2 x T8
    wire T54 = T2 & T8;
    // T55 = T41 x T39
    wire T55 = T41 & T39;
    // T56 = T55 + T54
    wire T56 = T55 ^ T54;
    // T57 = T16 x T14
    wire T57 = T16 & T14;
    // T58 = T57 + T54
    wire T58 = T57 ^ T54;
    // T59 = T46 + T45
    wire T59 = T46 ^ T45;
    // T60 = T48 + T42
    wire T60 = T48 ^ T42;
    // T61 = T51 + T50
    wire T61 = T51 ^ T50;
    // T62 = T53 + T58
    wire T62 = T53 ^ T58;
    // T63 = T59 + T56
    wire T63 = T59 ^ T56;
    // T64 = T60 + T58
    wire T64 = T60 ^ T58;
    // T65 = T61 + T56
    wire T65 = T61 ^ T56;
    // T66 = T62 + T43
    wire T66 = T62 ^ T43;
    // T67 = T65 + T66
    wire T67 = T65 ^ T66;
    // T68 = T65 x T63
    wire T68 = T65 & T63;
    // T69 = T64 + T68
    wire T69 = T64 ^ T68;
    // T70 = T63 + T64
    wire T70 = T63 ^ T64;
    // T71 = T66 + T68
    wire T71 = T66 ^ T68;
    // T72 = T71 x T70
    wire T72 = T71 & T70;
    // T73 = T69 x T67
    wire T73 = T69 & T67;
    // T74 = T63 x T66
    wire T74 = T63 & T66;
    // T75 = T70 x T74
    wire T75 = T70 & T74;
    // T76 = T70 + T68
    wire T76 = T70 ^ T68;
    // T77 = T64 x T65
    wire T77 = T64 & T65;
    // T78 = T67 x T77
    wire T78 = T67 & T77;
    // T79 = T67 + T68
    wire T79 = T67 ^ T68;
    // T80 = T64 + T72
    wire T80 = T64 ^ T72;
    // T81 = T75 + T76
    wire T81 = T75 ^ T76;
    // T82 = T66 + T73
    wire T82 = T66 ^ T73;
    // T83 = T78 + T79
    wire T83 = T78 ^ T79;
    // T84 = T81 + T83
    wire T84 = T81 ^ T83;
    // T85 = T80 + T82
    wire T85 = T80 ^ T82;
    // T86 = T80 + T81
    wire T86 = T80 ^ T81;
    // T87 = T82 + T83
    wire T87 = T82 ^ T83;
    // T88 = T85 + T84
    wire T88 = T85 ^ T84;
    // T89 = T87 x T5
    wire T89 = T87 & T5;
    // T90 = T83 x T11
    wire T90 = T83 & T11;
    // T91 = T82 x U7
    wire T91 = T82 & x[7];
    // T92 = T86 x T21
    wire T92 = T86 & T21;
    // T93 = T81 x T4
    wire T93 = T81 & T4;
    // T94 = T80 x T17
    wire T94 = T80 & T17;
    // T95 = T85 x T8
    wire T95 = T85 & T8;
    // T96 = T88 x T39
    wire T96 = T88 & T39;
    // T97 = T84 x T14
    wire T97 = T84 & T14;
    // T98 = T87 x T19
    wire T98 = T87 & T19;
    // T99 = T83 x T20
    wire T99 = T83 & T20;
    // T100 = T82 x T10
    wire T100 = T82 & T10;
    // T101 = T86 x T7
    wire T101 = T86 & T7;
    // T102 = T81 x T9
    wire T102 = T81 & T9;
    // T103 = T80 x T22
    wire T103 = T80 & T22;
    // T104 = T85 x T2
    wire T104 = T85 & T2;
    // T105 = T88 x T41
    wire T105 = T88 & T41;
    // T106 = T84 x T16
    wire T106 = T84 & T16;
    // T107 = T104 + T105
    wire T107 = T104 ^ T105;
    // T108 = T93 + T99
    wire T108 = T93 ^ T99;
    // T109 = T96 + T107
    wire T109 = T96 ^ T107;
    // T110 = T98 + T108
    wire T110 = T98 ^ T108;
    // T111 = T91 + T101
    wire T111 = T91 ^ T101;
    // T112 = T89 + T92
    wire T112 = T89 ^ T92;
    // T113 = T107 + T112
    wire T113 = T107 ^ T112;
    // T114 = T90 + T110
    wire T114 = T90 ^ T110;
    // T115 = T89 + T95
    wire T115 = T89 ^ T95;
    // T116 = T94 + T102
    wire T116 = T94 ^ T102;
    // T117 = T97 + T103
    wire T117 = T97 ^ T103;
    // T118 = T91 + T114
    wire T118 = T91 ^ T114;
    // T119 = T111 + T117
    wire T119 = T111 ^ T117;
    // T120 = T100 + T108
    wire T120 = T100 ^ T108;
    // T121 = T92 + T95
    wire T121 = T92 ^ T95;
    // T122 = T110 + T121
    wire T122 = T110 ^ T121;
    // T123 = T106 + T119
    wire T123 = T106 ^ T119;
    // T124 = T104 + T115
    wire T124 = T104 ^ T115;
    // T125 = T111 + T116
    wire T125 = T111 ^ T116;
    // S0 = T109 + T122
    wire S0 = T109 ^ T122;
    // S2 = T123 # T124
    wire S2 = T123 ^~ T124;
    // T128 = T94 + T107
    wire T128 = T94 ^ T107;
    // S3 = T113 + T114
    wire S3 = T113 ^ T114;
    // S4 = T118 + T128
    wire S4 = T118 ^ T128;
    // T131 = T93 + T101
    wire T131 = T93 ^ T101;
    // T132 = T112 + T120
    wire T132 = T112 ^ T120;
    // S7 = T113 # T125
    wire S7 = T113 ^~ T125;
    // T134 = T97 + T116
    wire T134 = T97 ^ T116;
    // T135 = T131 + T134
    wire T135 = T131 ^ T134;
    // T136 = T93 + T115
    wire T136 = T93 ^ T115;
    // S6 = T109 # T135
    wire S6 = T109 ^~ T135;
    // T138 = T119 + T132
    wire T138 = T119 ^ T132;
    // S5 = T109 + T138
    wire S5 = T109 ^ T138;
    // T140 = T114 + T136
    wire T140 = T114 ^ T136;
    // S1 = T109 # T140
    wire S1 = T109 ^~ T140;

    assign out = {S0, S1, S2, S3, S4, S5, S6, S7};
endmodule